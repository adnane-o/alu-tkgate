//: version "1.6f"
//: script "/home/xidus/mips/mips-single.gss"


module and6(I4, I3, I2, I1, Z, I5, I0);
//: interface  /sz:(87, 58) /bd:[ Ti0>I1(20/87) Ti1>I2(34/87) Ti2>I3(49/87) Ti3>I4(64/87) Ti4>I5(79/87) Ti5>I0(8/87) Bo0<Z(46/87) ]
input I2;    //: /sn:0 {0}(278,95)(278,165)(302,165)(302,175){1}
input I4;    //: /sn:0 {0}(381,95)(381,167)(406,167)(406,177){1}
input I1;    //: /sn:0 {0}(243,92)(243,131)(222,131)(222,174){1}
output Z;    //: /sn:0 /dp:1 {0}(305,287)(305,346){1}
input I5;    //: /sn:0 {0}(411,94)(411,177){1}
input I0;    //: /sn:0 {0}(217,92)(217,174){1}
input I3;    //: /sn:0 {0}(333,95)(333,165)(307,165)(307,175){1}
wire w8;    //: /sn:0 {0}(409,198)(409,257)(308,257)(308,266){1}
wire w2;    //: /sn:0 {0}(220,195)(220,256)(301,256)(301,266){1}
wire w5;    //: /sn:0 {0}(305,196)(305,266){1}
//: enddecls

  and g8 (.I0(I2), .I1(I3), .Z(w5));   //: @(305,186) /sn:0 /R:3 /w:[ 1 1 0 ]
  //: input g4 (I4) @(381,93) /sn:0 /R:3 /w:[ 0 ]
  //: input g3 (I3) @(333,93) /sn:0 /R:3 /w:[ 0 ]
  //: input g2 (I2) @(278,93) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (I1) @(243,90) /sn:0 /R:3 /w:[ 0 ]
  and g10 (.I0(w2), .I1(w5), .I2(w8), .Z(Z));   //: @(305,277) /sn:0 /R:3 /w:[ 1 1 1 0 ]
  //: output g6 (Z) @(305,343) /sn:0 /R:3 /w:[ 1 ]
  and g9 (.I0(I4), .I1(I5), .Z(w8));   //: @(409,188) /sn:0 /R:3 /w:[ 1 1 0 ]
  and g7 (.I0(I0), .I1(I1), .Z(w2));   //: @(220,185) /sn:0 /R:3 /w:[ 1 1 0 ]
  //: input g5 (I5) @(411,92) /sn:0 /R:3 /w:[ 0 ]
  //: input g0 (I0) @(217,90) /sn:0 /R:3 /w:[ 0 ]

endmodule

module imemory(MemData, Read, WriteData, Write, Addr);
//: interface  /sz:(89, 94) /bd:[ Ti0>Read(24/89) Ti1>Write(61/89) Li0>WriteData[31:0](76/94) Li1>Addr[31:0](27/94) Ro0<MemData[31:0](36/94) ]
supply0 w0;    //: /sn:0 {0}(240,191)(240,176){1}
input Read;    //: /sn:0 {0}(214,244)(254,244)(254,176){1}
input [31:0] Addr;    //: /sn:0 {0}(124,166)(167,166)(167,149){1}
//: {2}(167,148)(167,122){3}
input [31:0] WriteData;    //: /sn:0 {0}(327,75)(335,75)(335,128){1}
input Write;    //: /sn:0 {0}(201,50)(247,50)(247,91){1}
//: {2}(249,93)(350,93)(350,136)(340,136){3}
//: {4}(247,95)(247,126){5}
output [31:0] MemData;    //: /sn:0 {0}(335,144)(335,172){1}
//: {2}(337,174)(370,174){3}
//: {4}(333,174)(279,174)(279,149)(264,149){5}
wire [29:0] w5;    //: /sn:0 {0}(171,149)(229,149){1}
//: enddecls

  //: comment g4 /dolink:0 /link:"" @(160,98) /sn:0
  //: /line:"div4"
  //: /end
  //: output g8 (MemData) @(367,174) /sn:0 /w:[ 3 ]
  tran g3(.Z(w5), .I(Addr[31:2]));   //: @(165,149) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: supply0 g2 (w0) @(240,197) /sn:0 /w:[ 0 ]
  //: joint g11 (Write) @(247, 93) /w:[ 2 1 -1 4 ]
  //: joint g10 (MemData) @(335, 174) /w:[ 2 1 4 -1 ]
  //: input g6 (Read) @(212,244) /sn:0 /w:[ 0 ]
  ram m1 (.A(w5), .D(MemData), .WE(!Write), .OE(!Read), .CS(w0));   //: @(247,150) /sn:0 /w:[ 1 5 5 1 1 ]
  //: input g7 (WriteData) @(325,75) /sn:0 /w:[ 0 ]
  bufif1 g9 (.Z(MemData), .I(WriteData), .E(Write));   //: @(335,134) /sn:0 /R:3 /w:[ 0 1 3 ]
  //: input g5 (Write) @(199,50) /sn:0 /w:[ 0 ]
  //: input g0 (Addr) @(122,166) /sn:0 /w:[ 0 ]

endmodule

module dmemory(MemData, Read, WriteData, Write, Addr);
//: interface  /sz:(89, 94) /bd:[ Ti0>Read(24/89) Ti1>Write(61/89) Li0>WriteData[31:0](76/94) Li1>Addr[31:0](27/94) Ro0<MemData[31:0](36/94) ]
supply0 w0;    //: /sn:0 {0}(240,191)(240,176){1}
input Read;    //: /sn:0 {0}(214,244)(254,244)(254,176){1}
input [31:0] Addr;    //: /sn:0 {0}(124,166)(167,166)(167,149){1}
//: {2}(167,148)(167,122){3}
input [31:0] WriteData;    //: /sn:0 {0}(327,75)(335,75)(335,128){1}
input Write;    //: /sn:0 {0}(201,50)(247,50)(247,91){1}
//: {2}(249,93)(350,93)(350,136)(340,136){3}
//: {4}(247,95)(247,126){5}
output [31:0] MemData;    //: /sn:0 {0}(335,144)(335,172){1}
//: {2}(337,174)(370,174){3}
//: {4}(333,174)(279,174)(279,149)(264,149){5}
wire [29:0] w5;    //: /sn:0 {0}(171,149)(229,149){1}
//: enddecls

  //: comment g4 /dolink:0 /link:"" @(160,98) /sn:0
  //: /line:"div4"
  //: /end
  //: output g8 (MemData) @(367,174) /sn:0 /w:[ 3 ]
  tran g3(.Z(w5), .I(Addr[31:2]));   //: @(165,149) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: supply0 g2 (w0) @(240,197) /sn:0 /w:[ 0 ]
  //: joint g11 (Write) @(247, 93) /w:[ 2 1 -1 4 ]
  //: joint g10 (MemData) @(335, 174) /w:[ 2 1 4 -1 ]
  ram m1 (.A(w5), .D(MemData), .WE(!Write), .OE(!Read), .CS(w0));   //: @(247,150) /sn:0 /w:[ 1 5 5 1 1 ]
  //: input g6 (Read) @(212,244) /sn:0 /w:[ 0 ]
  //: input g7 (WriteData) @(325,75) /sn:0 /w:[ 0 ]
  bufif1 g9 (.Z(MemData), .I(WriteData), .E(Write));   //: @(335,134) /sn:0 /R:3 /w:[ 0 1 3 ]
  //: input g5 (Write) @(199,50) /sn:0 /w:[ 0 ]
  //: input g0 (Addr) @(122,166) /sn:0 /w:[ 0 ]

endmodule

module ALU(Z, B, zero, ALUOp, A);
//: interface  /sz:(83, 90) /bd:[ Li0>B[31:0](55/90) Li1>A[31:0](18/90) Bi0>ALUOp[2:0](38/83) Ro0<Z[31:0](41/90) Ro1<zero(6/90) ]
input [31:0] B;    //: /sn:0 {0}(78,97)(153,97){1}
//: {2}(157,97)(271,97){3}
//: {4}(275,97)(295,97)(295,187){5}
//: {6}(273,99)(273,187){7}
//: {8}(155,99)(155,125){9}
input [31:0] A;    //: /sn:0 {0}(89,82)(124,82){1}
//: {2}(128,82)(266,82){3}
//: {4}(270,82)(290,82)(290,187){5}
//: {6}(268,84)(268,187){7}
//: {8}(126,84)(126,168){9}
supply0 [30:0] w3;    //: /sn:0 {0}(446,279)(446,272)(389,272){1}
output zero;    //: /sn:0 /dp:1 {0}(243,378)(295,378){1}
output [31:0] Z;    //: /sn:0 /dp:1 {0}(310,313)(310,343)(347,343){1}
input [2:0] ALUOp;    //: /sn:0 {0}(192,300)(237,300){1}
//: {2}(238,300)(287,300){3}
supply0 [31:0] w10;    //: /sn:0 {0}(372,232)(372,222)(357,222)(357,259)(321,259){1}
//: {2}(317,259)(306,259)(306,267){3}
//: {4}(308,269)(313,269)(313,284){5}
//: {6}(306,271)(306,284){7}
//: {8}(319,261)(319,284){9}
wire w14;    //: /sn:0 {0}(238,295)(238,182)(214,182){1}
//: {2}(212,180)(212,115)(160,115)(160,125){3}
//: {4}(210,182)(166,182){5}
wire [31:0] w16;    //: /sn:0 {0}(271,208)(271,269)(286,269)(286,284){1}
wire w15;    //: /sn:0 {0}(118,182)(108,182){1}
wire [31:0] w19;    //: /sn:0 {0}(293,208)(293,284){1}
wire w0;    //: /sn:0 {0}(330,250)(406,250)(406,282)(389,282){1}
wire [31:0] w8;    //: /sn:0 {0}(158,146)(158,168){1}
wire [31:0] w2;    //: /sn:0 {0}(383,277)(333,277)(333,284){1}
wire [31:0] w13;    //: /sn:0 {0}(142,197)(142,242){1}
//: {2}(144,244)(297,244){3}
//: {4}(301,244)(326,244)(326,249){5}
//: {6}(326,250)(326,284){7}
//: {8}(299,246)(299,284){9}
//: {10}(142,246)(142,378)(222,378){11}
//: enddecls

  //: supply0 g4 (w10) @(372,238) /sn:0 /w:[ 0 ]
  and g8 (.I0(A), .I1(B), .Z(w16));   //: @(271,198) /sn:0 /R:3 /w:[ 7 7 0 ]
  mux g3 (.I0(w16), .I1(w19), .I2(w13), .I3(w10), .I4(w10), .I5(w10), .I6(w13), .I7(w2), .S(ALUOp), .Z(Z));   //: @(310,300) /sn:0 /w:[ 1 1 9 7 5 9 7 1 3 0 ]
  xor g13 (.I0(B), .I1(w14), .Z(w8));   //: @(158,136) /sn:0 /R:3 /w:[ 9 3 0 ]
  //: output g2 (Z) @(344,343) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(76,97) /sn:0 /w:[ 0 ]
  //: joint g11 (B) @(273, 97) /w:[ 4 -1 3 6 ]
  //: joint g16 (w13) @(299, 244) /w:[ 4 -1 3 8 ]
  //: joint g10 (A) @(268, 82) /w:[ 4 -1 3 6 ]
  //: output g19 (zero) @(292,378) /sn:0 /w:[ 1 ]
  //: input g6 (ALUOp) @(190,300) /sn:0 /w:[ 0 ]
  tran g7(.Z(w14), .I(ALUOp[2]));   //: @(238,298) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  or g9 (.I0(A), .I1(B), .Z(w19));   //: @(293,198) /sn:0 /R:3 /w:[ 5 5 0 ]
  //: joint g15 (w14) @(212, 182) /w:[ 1 2 4 -1 ]
  nor g20 (.I0(w13), .Z(zero));   //: @(233,378) /sn:0 /w:[ 11 0 ]
  //: joint g17 (w10) @(306, 269) /w:[ 4 3 -1 6 ]
  add g5 (.A(A), .B(w8), .S(w13), .CI(w14), .CO(w15));   //: @(142,184) /sn:0 /w:[ 9 1 0 5 0 ]
  //: joint g14 (B) @(155, 97) /w:[ 2 -1 1 8 ]
  //: joint g21 (w13) @(142, 244) /w:[ 2 1 -1 10 ]
  tran g24(.Z(w0), .I(w13[31]));   //: @(324,250) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  //: supply0 g23 (w3) @(446,285) /sn:0 /w:[ 0 ]
  //: input g0 (A) @(87,82) /sn:0 /w:[ 0 ]
  concat g22 (.I0(w0), .I1(w3), .Z(w2));   //: @(384,277) /sn:0 /R:2 /w:[ 1 1 0 ] /dr:1
  //: joint g12 (A) @(126, 82) /w:[ 2 -1 1 8 ]
  //: joint g18 (w10) @(319, 259) /w:[ 1 -1 2 8 ]

endmodule

module control(RegWrite, MemToReg, ALUSrc, RegDest, ALUOp, Branch, MemWrite, MemRead, Op);
//: interface  /sz:(111, 110) /bd:[ Bi0>Op[5:0](62/111) Lo0<Branch(27/110) Ro0<RegDest(6/110) Ro1<MemRead(26/110) Ro2<MemToReg(16/110) Ro3<MemWrite(37/110) Ro4<ALUOp[1:0](65/110) Ro5<ALUSrc(80/110) Ro6<RegWrite(92/110) ]
output MemToReg;    //: /sn:0 {0}(301,459)(271,459)(271,412){1}
//: {2}(273,410)(598,410){3}
//: {4}(271,408)(271,324){5}
output RegDest;    //: /sn:0 {0}(552,532)(153,532)(153,387){1}
//: {2}(155,385)(529,385){3}
//: {4}(153,383)(153,364){5}
//: {6}(155,362)(600,362){7}
//: {8}(153,360)(153,324){9}
output MemWrite;    //: /sn:0 {0}(599,482)(393,482)(393,437){1}
//: {2}(395,435)(530,435){3}
//: {4}(393,433)(393,324){5}
output Branch;    //: /sn:0 {0}(530,440)(512,440){1}
//: {2}(510,438)(510,382){3}
//: {4}(512,380)(529,380){5}
//: {6}(510,378)(510,326){7}
//: {8}(510,442)(510,507){9}
//: {10}(512,509)(599,509){11}
//: {12}(510,511)(510,542)(552,542){13}
output ALUSrc;    //: /sn:0 {0}(599,383)(550,383){1}
input [5:0] Op;    //: /sn:0 {0}(38,60)(64,60)(64,65){1}
//: {2}(64,66)(64,81){3}
//: {4}(64,82)(64,97){5}
//: {6}(64,98)(64,113){7}
//: {8}(64,114)(64,129){9}
//: {10}(64,130)(64,144){11}
//: {12}(64,145)(64,167){13}
output [1:0] ALUOp;    //: /sn:0 /dp:1 {0}(558,537)(598,537){1}
output RegWrite;    //: /sn:0 /dp:1 {0}(551,438)(600,438){1}
output MemRead;    //: /sn:0 /dp:1 {0}(317,459)(600,459){1}
wire w6;    //: /sn:0 {0}(355,264)(355,68){1}
//: {2}(357,66)(472,66)(472,204){3}
//: {4}(353,66)(235,66){5}
//: {6}(231,66)(117,66){7}
//: {8}(113,66)(68,66){9}
//: {10}(115,68)(115,204){11}
//: {12}(233,68)(233,264){13}
wire w45;    //: /sn:0 {0}(396,220)(396,264){1}
wire w4;    //: /sn:0 {0}(411,264)(411,132){1}
//: {2}(413,130)(528,130)(528,204){3}
//: {4}(409,130)(291,130){5}
//: {6}(287,130)(173,130){7}
//: {8}(169,130)(68,130){9}
//: {10}(171,132)(171,204){11}
//: {12}(289,132)(289,264){13}
wire w51;    //: /sn:0 {0}(528,220)(528,266){1}
wire w3;    //: /sn:0 {0}(68,114)(154,114){1}
//: {2}(158,114)(272,114){3}
//: {4}(276,114)(394,114){5}
//: {6}(398,114)(513,114)(513,266){7}
//: {8}(396,116)(396,204){9}
//: {10}(274,116)(274,204){11}
//: {12}(156,116)(156,204){13}
wire w37;    //: /sn:0 {0}(245,220)(245,264){1}
wire w43;    //: /sn:0 {0}(367,220)(367,264){1}
wire w31;    //: /sn:0 {0}(141,220)(141,264){1}
wire w41;    //: /sn:0 {0}(274,220)(274,264){1}
wire w8;    //: /sn:0 {0}(186,220)(186,264){1}
wire w35;    //: /sn:0 {0}(171,220)(171,264){1}
wire w53;    //: /sn:0 {0}(543,220)(543,266){1}
wire w49;    //: /sn:0 {0}(498,220)(498,266){1}
wire w2;    //: /sn:0 /dp:1 {0}(381,264)(381,100){1}
//: {2}(383,98)(498,98)(498,204){3}
//: {4}(379,98)(261,98){5}
//: {6}(257,98)(143,98){7}
//: {8}(139,98)(68,98){9}
//: {10}(141,100)(141,204){11}
//: {12}(259,100)(259,204){13}
wire w10;    //: /sn:0 {0}(484,220)(484,266){1}
wire w33;    //: /sn:0 {0}(156,220)(156,264){1}
wire w5;    //: /sn:0 {0}(426,264)(426,147){1}
//: {2}(428,145)(543,145)(543,204){3}
//: {4}(424,145)(306,145){5}
//: {6}(302,145)(188,145){7}
//: {8}(184,145)(68,145){9}
//: {10}(186,147)(186,204){11}
//: {12}(304,147)(304,264){13}
wire w47;    //: /sn:0 {0}(472,220)(472,266){1}
wire w29;    //: /sn:0 {0}(127,220)(127,264){1}
wire w9;    //: /sn:0 {0}(484,204)(484,82)(369,82){1}
//: {2}(365,82)(247,82){3}
//: {4}(243,82)(129,82){5}
//: {6}(125,82)(68,82){7}
//: {8}(127,84)(127,204){9}
//: {10}(245,84)(245,204){11}
//: {12}(367,84)(367,204){13}
wire w39;    //: /sn:0 {0}(259,220)(259,264){1}
wire w26;    //: /sn:0 {0}(115,220)(115,264){1}
//: enddecls

  //: output g4 (RegWrite) @(597,438) /sn:0 /w:[ 1 ]
  tran g8(.Z(w3), .I(Op[2]));   //: @(62,114) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  //: joint g51 (Branch) @(510, 380) /w:[ 4 6 -1 3 ]
  buf g55 (.I(MemToReg), .Z(MemRead));   //: @(307,459) /sn:0 /w:[ 0 0 ]
  //: output g3 (MemToReg) @(595,410) /sn:0 /w:[ 3 ]
  //: joint g37 (w2) @(259, 98) /w:[ 5 -1 6 12 ]
  //: joint g34 (w4) @(171, 130) /w:[ 7 -1 8 10 ]
  not g13 (.I(w2), .Z(w31));   //: @(141,210) /sn:0 /R:3 /w:[ 11 0 ]
  //: output g2 (ALUSrc) @(596,383) /sn:0 /w:[ 0 ]
  //: joint g59 (Branch) @(510, 509) /w:[ 10 9 -1 12 ]
  //: output g1 (RegDest) @(597,362) /sn:0 /w:[ 7 ]
  not g16 (.I(w9), .Z(w37));   //: @(245,210) /sn:0 /R:3 /w:[ 11 0 ]
  not g11 (.I(w6), .Z(w26));   //: @(115,210) /sn:0 /R:3 /w:[ 11 0 ]
  and g50 (.I0(!Branch), .I1(!RegDest), .Z(ALUSrc));   //: @(540,383) /sn:0 /w:[ 5 3 1 ]
  not g28 (.I(w5), .Z(w8));   //: @(186,210) /sn:0 /R:3 /w:[ 11 0 ]
  tran g10(.Z(w5), .I(Op[0]));   //: @(62,145) /sn:0 /R:2 /w:[ 9 12 11 ] /ss:1
  //: joint g32 (w2) @(141, 98) /w:[ 7 -1 8 10 ]
  not g27 (.I(w5), .Z(w53));   //: @(543,210) /sn:0 /R:3 /w:[ 3 0 ]
  not g19 (.I(w3), .Z(w41));   //: @(274,210) /sn:0 /R:3 /w:[ 11 0 ]
  and6 rform (.I0(w26), .I5(w8), .I4(w35), .I3(w33), .I2(w31), .I1(w29), .Z(RegDest));   //: @(107, 265) /sz:(87, 58) /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Bo0<9 ]
  and6 sw (.I0(w6), .I5(w5), .I4(w4), .I3(w45), .I2(w2), .I1(w43), .Z(MemWrite));   //: @(347, 265) /sz:(87, 58) /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>1 Ti4>0 Ti5>1 Bo0<5 ]
  //: joint g38 (w3) @(274, 114) /w:[ 4 -1 3 10 ]
  tran g6(.Z(w9), .I(Op[4]));   //: @(62,82) /sn:0 /R:2 /w:[ 7 4 3 ] /ss:1
  //: joint g57 (RegDest) @(153, 385) /w:[ 2 4 -1 1 ]
  //: joint g53 (MemToReg) @(271, 410) /w:[ 2 4 -1 1 ]
  tran g9(.Z(w4), .I(Op[1]));   //: @(62,130) /sn:0 /R:2 /w:[ 9 10 9 ] /ss:1
  tran g7(.Z(w2), .I(Op[3]));   //: @(62,98) /sn:0 /R:2 /w:[ 9 6 5 ] /ss:1
  //: joint g31 (w9) @(127, 82) /w:[ 5 -1 6 8 ]
  not g20 (.I(w9), .Z(w43));   //: @(367,210) /sn:0 /R:3 /w:[ 13 0 ]
  not g15 (.I(w4), .Z(w35));   //: @(171,210) /sn:0 /R:3 /w:[ 11 0 ]
  and6 lw (.I0(w6), .I5(w5), .I4(w4), .I3(w41), .I2(w39), .I1(w37), .Z(MemToReg));   //: @(225, 265) /sz:(87, 58) /p:[ Ti0>13 Ti1>13 Ti2>13 Ti3>1 Ti4>1 Ti5>1 Bo0<5 ]
  //: joint g39 (w9) @(367, 82) /w:[ 1 -1 2 12 ]
  //: output g48 (ALUOp) @(595,537) /sn:0 /w:[ 1 ]
  //: joint g43 (w4) @(411, 130) /w:[ 2 -1 4 1 ]
  not g29 (.I(w9), .Z(w10));   //: @(484,210) /sn:0 /R:3 /w:[ 0 0 ]
  not g25 (.I(w2), .Z(w49));   //: @(498,210) /sn:0 /R:3 /w:[ 3 0 ]
  //: joint g17 (w6) @(233, 66) /w:[ 5 -1 6 12 ]
  and g52 (.I0(!MemWrite), .I1(!Branch), .Z(RegWrite));   //: @(541,438) /sn:0 /w:[ 3 0 0 ]
  //: joint g42 (w2) @(381, 98) /w:[ 2 -1 4 1 ]
  //: joint g56 (MemWrite) @(393, 435) /w:[ 2 4 -1 1 ]
  not g14 (.I(w3), .Z(w33));   //: @(156,210) /sn:0 /R:3 /w:[ 13 0 ]
  tran g5(.Z(w6), .I(Op[5]));   //: @(62,66) /sn:0 /R:2 /w:[ 9 2 1 ] /ss:1
  //: output g47 (Branch) @(596,509) /sn:0 /w:[ 11 ]
  //: joint g44 (w5) @(426, 145) /w:[ 2 -1 4 1 ]
  //: joint g36 (w9) @(245, 82) /w:[ 3 -1 4 10 ]
  not g24 (.I(w6), .Z(w47));   //: @(472,210) /sn:0 /R:3 /w:[ 3 0 ]
  //: joint g21 (w4) @(289, 130) /w:[ 5 -1 6 12 ]
  //: joint g41 (w6) @(355, 66) /w:[ 2 -1 4 1 ]
  not g23 (.I(w3), .Z(w45));   //: @(396,210) /sn:0 /R:3 /w:[ 9 0 ]
  //: joint g60 (Branch) @(510, 440) /w:[ 1 2 -1 8 ]
  //: joint g54 (RegDest) @(153, 362) /w:[ 6 8 -1 5 ]
  //: joint g40 (w3) @(396, 114) /w:[ 6 -1 5 8 ]
  //: output g46 (MemWrite) @(596,482) /sn:0 /w:[ 0 ]
  //: output g45 (MemRead) @(597,459) /sn:0 /w:[ 1 ]
  //: joint g35 (w5) @(186, 145) /w:[ 7 -1 8 10 ]
  not g26 (.I(w4), .Z(w51));   //: @(528,210) /sn:0 /R:3 /w:[ 3 0 ]
  //: joint g22 (w5) @(304, 145) /w:[ 5 -1 6 12 ]
  //: input g0 (Op) @(36,60) /sn:0 /w:[ 0 ]
  not g18 (.I(w2), .Z(w39));   //: @(259,210) /sn:0 /R:3 /w:[ 13 0 ]
  not g12 (.I(w9), .Z(w29));   //: @(127,210) /sn:0 /R:3 /w:[ 9 0 ]
  and6 beq (.I0(w47), .I5(w53), .I4(w51), .I3(w3), .I2(w49), .I1(w10), .Z(Branch));   //: @(464, 267) /sz:(87, 58) /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>7 Ti4>1 Ti5>1 Bo0<7 ]
  //: joint g33 (w3) @(156, 114) /w:[ 2 -1 1 12 ]
  //: joint g30 (w6) @(115, 66) /w:[ 7 -1 8 10 ]
  concat g49 (.I0(Branch), .I1(RegDest), .Z(ALUOp));   //: @(557,537) /sn:0 /w:[ 13 0 0 ] /dr:0

endmodule

module reg4(CLK, SB, WEN, SA, DA, ENA, CLR, WD, DB, WA, ENB);
//: interface  /sz:(102, 109) /bd:[ Ti0>WD[31:0](49/102) Li0>CLK(101/109) Li1>CLR(91/109) Li2>WEN(72/109) Li3>WA[1:0](61/109) Li4>ENB(46/109) Li5>ENA(35/109) Li6>SB[1:0](21/109) Li7>SA[1:0](9/109) Bo0<DB[31:0](78/102) Bo1<DA[31:0](30/102) ]
input ENB;    //: /sn:0 {0}(573,526)(537,526)(537,563){1}
input [1:0] WA;    //: /sn:0 {0}(36,377)(78,377){1}
input [31:0] WD;    //: /sn:0 {0}(84,109)(215,109){1}
//: {2}(219,109)(379,109){3}
//: {4}(383,109)(532,109){5}
//: {6}(536,109)(673,109)(673,212){7}
//: {8}(534,111)(534,212){9}
//: {10}(381,111)(381,212){11}
//: {12}(217,111)(217,212){13}
input [1:0] SB;    //: /sn:0 {0}(444,502)(483,502){1}
input CLR;    //: /sn:0 {0}(43,304)(271,304){1}
//: {2}(275,304)(437,304){3}
//: {4}(441,304)(589,304){5}
//: {6}(593,304)(731,304)(731,217)(712,217){7}
//: {8}(591,302)(591,217)(573,217){9}
//: {10}(439,302)(439,217)(420,217){11}
//: {12}(273,302)(273,217)(256,217){13}
input [1:0] SA;    //: /sn:0 {0}(194,502)(255,502){1}
input WEN;    //: /sn:0 {0}(34,340)(91,340)(91,353){1}
output [31:0] DB;    //: /sn:0 {0}(585,568)(545,568){1}
input CLK;    //: /sn:0 {0}(43,283)(167,283){1}
//: {2}(171,283)(328,283){3}
//: {4}(332,283)(485,283){5}
//: {6}(489,283)(627,283)(627,222)(636,222){7}
//: {8}(487,281)(487,222)(497,222){9}
//: {10}(330,281)(330,222)(344,222){11}
//: {12}(169,281)(169,222)(180,222){13}
output [31:0] DA;    //: /sn:0 /dp:1 {0}(309,572)(344,572){1}
input ENA;    //: /sn:0 {0}(332,528)(301,528)(301,567){1}
wire w14;    //: /sn:0 {0}(107,395)(722,395)(722,227)(712,227){1}
wire [31:0] w15;    //: /sn:0 {0}(673,233)(673,457)(526,457){1}
//: {2}(522,457)(296,457)(296,486){3}
//: {4}(524,459)(524,471)(524,471)(524,486){5}
wire [31:0] w0;    //: /sn:0 {0}(217,233)(217,431)(258,431){1}
//: {2}(262,431)(488,431)(488,486){3}
//: {4}(260,433)(260,460)(260,460)(260,486){5}
wire [31:0] w23;    //: /sn:0 {0}(278,515)(278,572)(293,572){1}
wire w8;    //: /sn:0 {0}(107,359)(265,359)(265,227)(256,227){1}
wire [31:0] w10;    //: /sn:0 {0}(534,233)(534,447)(514,447){1}
//: {2}(510,447)(284,447)(284,486){3}
//: {4}(512,449)(512,466)(512,466)(512,486){5}
wire [31:0] w27;    //: /sn:0 {0}(506,515)(506,568)(529,568){1}
wire w13;    //: /sn:0 {0}(107,383)(585,383)(585,227)(573,227){1}
wire [31:0] w5;    //: /sn:0 {0}(381,233)(381,436){1}
//: {2}(383,438)(500,438)(500,486){3}
//: {4}(379,438)(272,438)(272,486){5}
wire w9;    //: /sn:0 {0}(107,371)(430,371)(430,227)(420,227){1}
//: enddecls

  mux g4 (.I0(w0), .I1(w5), .I2(w10), .I3(w15), .S(SA), .Z(w23));   //: @(278,502) /sn:0 /w:[ 5 5 3 3 1 0 ]
  //: joint g8 (w10) @(512, 447) /w:[ 1 -1 2 4 ]
  register g3 (.Q(w15), .D(WD), .EN(!w14), .CLR(!CLR), .CK(CLK));   //: @(673,222) /sn:0 /w:[ 0 7 1 7 7 ]
  //: joint g13 (CLK) @(487, 283) /w:[ 6 8 5 -1 ]
  register g2 (.Q(w10), .D(WD), .EN(!w13), .CLR(!CLR), .CK(CLK));   //: @(534,222) /sn:0 /w:[ 0 9 1 9 9 ]
  register g1 (.Q(w5), .D(WD), .EN(!w9), .CLR(!CLR), .CK(CLK));   //: @(381,222) /sn:0 /w:[ 0 11 1 11 11 ]
  //: joint g11 (CLK) @(169, 283) /w:[ 2 12 1 -1 ]
  //: joint g16 (CLR) @(439, 304) /w:[ 4 10 3 -1 ]
  //: input g10 (CLK) @(41,283) /sn:0 /w:[ 0 ]
  bufif1 g28 (.Z(DA), .I(w23), .E(ENA));   //: @(299,572) /sn:0 /w:[ 0 1 1 ]
  demux g19 (.I(WA), .E(WEN), .Z0(w8), .Z1(w9), .Z2(w13), .Z3(w14));   //: @(91,377) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 ]
  bufif1 g27 (.Z(DB), .I(w27), .E(ENB));   //: @(535,568) /sn:0 /w:[ 1 1 1 ]
  //: input g32 (SB) @(442,502) /sn:0 /w:[ 0 ]
  //: joint g6 (w0) @(260, 431) /w:[ 2 -1 1 4 ]
  //: joint g7 (w5) @(381, 438) /w:[ 2 1 4 -1 ]
  //: joint g9 (w15) @(524, 457) /w:[ 1 -1 2 4 ]
  //: joint g15 (CLR) @(273, 304) /w:[ 2 12 1 -1 ]
  //: input g20 (WEN) @(32,340) /sn:0 /w:[ 0 ]
  //: input g31 (SA) @(192,502) /sn:0 /w:[ 0 ]
  //: joint g17 (CLR) @(591, 304) /w:[ 6 8 5 -1 ]
  //: output g25 (DA) @(341,572) /sn:0 /w:[ 1 ]
  //: input g29 (ENA) @(334,528) /sn:0 /R:2 /w:[ 0 ]
  mux g5 (.I0(w0), .I1(w5), .I2(w10), .I3(w15), .S(SB), .Z(w27));   //: @(506,502) /sn:0 /w:[ 3 3 5 5 1 0 ]
  //: input g14 (CLR) @(41,304) /sn:0 /w:[ 0 ]
  //: input g21 (WD) @(82,109) /sn:0 /w:[ 0 ]
  //: joint g24 (WD) @(534, 109) /w:[ 6 -1 5 8 ]
  //: joint g23 (WD) @(381, 109) /w:[ 4 -1 3 10 ]
  register g0 (.Q(w0), .D(WD), .EN(!w8), .CLR(!CLR), .CK(CLK));   //: @(217,222) /sn:0 /w:[ 0 13 1 13 13 ]
  //: joint g22 (WD) @(217, 109) /w:[ 2 -1 1 12 ]
  //: output g26 (DB) @(582,568) /sn:0 /w:[ 0 ]
  //: joint g12 (CLK) @(330, 283) /w:[ 4 10 3 -1 ]
  //: input g18 (WA) @(34,377) /sn:0 /w:[ 0 ]
  //: input g30 (ENB) @(575,526) /sn:0 /R:2 /w:[ 0 ]

endmodule

module main;    //: root_module
supply1 w4;    //: /sn:0 {0}(184,120)(169,120){1}
//: {2}(165,120)(150,120)(150,115){3}
//: {4}(167,122)(167,130)(184,130){5}
supply0 [31:0] w0;    //: /sn:0 {0}(-194,184)(-194,173)(-183,173){1}
supply0 w3;    //: /sn:0 /dp:1 {0}(-138,76)(-138,66)(-121,66)(-121,96){1}
supply0 w36;    //: /sn:0 {0}(-413,81)(-413,76)(-432,76)(-432,90){1}
supply1 [15:0] w25;    //: /sn:0 {0}(99,248)(99,261)(108,261){1}
supply0 w11;    //: /sn:0 /dp:1 {0}(-41,95)(-41,85)(-26,85)(-26,95){1}
supply1 w5;    //: /sn:0 {0}(-158,54)(-158,96){1}
supply0 w9;    //: /sn:0 {0}(-243,83)(-243,78)(-271,78)(-271,86){1}
supply0 w42;    //: /sn:0 {0}(-194,322)(-194,312)(-210,312)(-210,334){1}
wire [31:0] w6;    //: /sn:0 {0}(-507,92)(-507,98)(-446,98){1}
wire w7;    //: /sn:0 /dp:1 {0}(646,90)(646,-57)(80,-57){1}
wire w45;    //: /sn:0 {0}(-432,138)(-432,148){1}
wire [31:0] B;    //: /sn:0 /dp:1 {0}(307,259)(346,259)(346,277)(386,277){1}
wire [4:0] WA;    //: /sn:0 /dp:1 {0}(133,145)(184,145){1}
wire [31:0] w46;    //: /sn:0 /dp:1 {0}(-358,134)(-370,134)(-370,276)(-183,276)(-183,358)(-195,358){1}
wire [1:0] w60;    //: /sn:0 /dp:1 {0}(80,-29)(319,-29)(319,310)(239,310)(239,326){1}
wire w61;    //: /sn:0 {0}(80,-14)(294,-14)(294,236){1}
wire [31:0] IR;    //: /sn:0 /dp:1 {0}(-36,133)(4,133){1}
//: {2}(5,133)(23,133)(23,107)(41,107){3}
wire [31:0] nextPC;    //: /sn:0 {0}(-329,124)(-287,124){1}
wire w56;    //: /sn:0 {0}(-33,-67)(-381,-67)(-381,33)(-371,33){1}
wire [31:0] PC;    //: /sn:0 /dp:4 {0}(-224,374)(-242,374)(-242,186){1}
//: {2}(-242,182)(-242,126){3}
//: {4}(-240,124)(-183,124){5}
//: {6}(-244,124)(-266,124){7}
//: {8}(-244,184)(-466,184)(-466,130)(-446,130){9}
wire [15:0] w38;    //: /sn:0 {0}(129,264)(193,264){1}
wire [31:0] A;    //: /sn:0 /dp:1 {0}(218,197)(218,221)(350,221)(350,240)(386,240){1}
wire zero;    //: /sn:0 /dp:1 {0}(-371,38)(-392,38)(-392,435)(491,435)(491,228)(471,228){1}
wire w37;    //: /sn:0 {0}(92,269)(92,266)(108,266){1}
wire [31:0] Z;    //: /sn:0 /dp:1 {0}(471,263)(535,263)(535,163){1}
//: {2}(537,161)(582,161){3}
//: {4}(535,159)(535,75)(562,75){5}
wire w63;    //: /sn:0 /dp:1 {0}(-342,101)(-342,36)(-350,36){1}
wire [31:0] w21;    //: /sn:0 {0}(673,170)(683,170)(683,124)(548,124)(548,95)(562,95){1}
wire [31:0] WD;    //: /sn:0 /dp:1 {0}(591,85)(601,85)(601,46)(232,46)(232,82){1}
wire w58;    //: /sn:0 {0}(80,-78)(578,-78)(578,62){1}
wire [5:0] Inst;    //: /sn:0 /dp:1 {0}(47,132)(64,132)(64,375)(204,375){1}
wire [4:0] w28;    //: /sn:0 {0}(47,112)(83,112)(83,155)(104,155){1}
wire [4:0] SB;    //: /sn:0 {0}(184,102)(94,102){1}
//: {2}(90,102)(47,102){3}
//: {4}(92,104)(92,135)(104,135){5}
wire [31:0] w20;    //: /sn:0 {0}(582,210)(257,210){1}
//: {2}(255,208)(255,197){3}
//: {4}(255,212)(255,249)(278,249){5}
wire [31:0] w24;    //: /sn:0 {0}(199,269)(225,269){1}
//: {2}(229,269)(278,269){3}
//: {4}(227,271)(227,300)(-289,300)(-289,342)(-279,342){5}
wire [31:0] w1;    //: /sn:0 {0}(-417,114)(-358,114){1}
wire [4:0] SA;    //: /sn:0 {0}(184,92)(47,92){1}
wire WEN;    //: /sn:0 /dp:1 {0}(80,-2)(140,-2)(140,156)(184,156){1}
wire [31:0] w30;    //: /sn:0 {0}(-92,133)(-57,133){1}
wire [15:0] w22;    //: /sn:0 {0}(5,137)(5,274)(91,274){1}
//: {2}(92,274)(193,274){3}
wire [5:0] Op;    //: /sn:0 /dp:1 {0}(47,82)(57,82)(57,47)(30,47)(30,17){1}
wire w12;    //: /sn:0 /dp:1 {0}(644,133)(644,111){1}
wire clk;    //: /sn:0 {0}(-342,-1)(-294,-1){1}
//: {2}(-290,-1)(-60,-1)(-60,183)(-48,183){3}
//: {4}(-44,183)(152,183){5}
//: {6}(156,183)(184,183){7}
//: {8}(154,185)(154,216)(513,216)(513,36)(641,36)(641,90){9}
//: {10}(-46,181)(-46,171){11}
//: {12}(-292,1)(-292,174)(-276,174)(-276,162){13}
wire [31:0] w49;    //: /sn:0 /dp:1 {0}(-224,342)(-258,342){1}
wire w57;    //: /sn:0 /dp:1 {0}(80,-68)(607,-68)(607,133){1}
wire [4:0] w44;    //: /sn:0 /dp:1 {0}(-295,414)(-268,414)(-268,380){1}
wire [2:0] ALUOp;    //: /sn:0 /dp:1 {0}(295,341)(425,341)(425,313){1}
wire [4:0] w13;    //: /sn:0 {0}(57,122)(47,122){1}
wire w48;    //: /sn:0 {0}(-210,382)(-210,392){1}
wire reset;    //: /sn:0 /dp:3 {0}(184,173)(16,173)(16,49)(-49,49){1}
//: {2}(-51,47)(-51,-33)(-279,-33){3}
//: {4}(-283,-33)(-339,-33){5}
//: {6}(-281,-31)(-281,86){7}
//: {8}(-51,51)(-51,95){9}
wire w50;    //: /sn:0 {0}(80,-88)(120,-88)(120,122){1}
//: enddecls

  and g8 (.I0(w25), .I1(w37), .Z(w38));   //: @(119,264) /sn:0 /w:[ 1 1 0 ]
  mux g4 (.I0(w20), .I1(w24), .S(w61), .Z(B));   //: @(294,259) /sn:0 /R:1 /w:[ 5 3 1 0 ]
  //: joint g37 (clk) @(-292, -1) /w:[ 2 -1 1 12 ]
  //: supply0 g34 (w3) @(-138,82) /sn:0 /w:[ 0 ]
  mux g13 (.I0(Z), .I1(w21), .S(w58), .Z(WD));   //: @(578,85) /sn:0 /R:1 /w:[ 5 1 1 0 ]
  concat g3 (.I0(w22), .I1(w38), .Z(w24));   //: @(198,269) /sn:0 /w:[ 3 1 0 ] /dr:0
  register IR (.Q(IR), .D(w30), .EN(w11), .CLR(!reset), .CK(clk));   //: @(-46,133) /R:1 /w:[ 0 1 0 9 11 ]
  and g2 (.I0(!clk), .I1(w7), .Z(w12));   //: @(644,101) /sn:0 /R:3 /w:[ 9 0 1 ]
  imemory imemory (.Read(w5), .Write(w3), .WriteData(w0), .Addr(PC), .MemData(w30));   //: @(-182, 97) /sz:(89, 94) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Li1>5 Ro0<0 ]
  register PC (.Q(PC), .D(nextPC), .EN(w9), .CLR(!reset), .CK(clk));   //: @(-276,124) /R:1 /w:[ 7 1 1 7 13 ]
  ALU g1 (.B(B), .A(A), .ALUOp(ALUOp), .Z(Z), .zero(zero));   //: @(387, 223) /sz:(83, 89) /sn:0 /p:[ Li0>1 Li1>1 Bi0>1 Ro0<0 Ro1<1 ]
  dmemory dmemory (.Read(w57), .Write(w12), .WriteData(w20), .Addr(Z), .MemData(w21));   //: @(583, 134) /sz:(89, 94) /sn:0 /p:[ Ti0>1 Ti1>0 Li0>0 Li1>3 Ro0<0 ]
  //: joint g11 (w4) @(167, 120) /w:[ 1 -1 2 4 ]
  add g16 (.A(PC), .B(w6), .S(w1), .CI(w36), .CO(w45));   //: @(-430,114) /sn:0 /R:1 /w:[ 9 1 0 1 0 ]
  //: supply1 g10 (w4) @(161,115) /sn:0 /w:[ 3 ]
  mux g28 (.I0(SB), .I1(w28), .S(w50), .Z(WA));   //: @(120,145) /sn:0 /R:1 /w:[ 5 1 1 0 ]
  //: joint g27 (PC) @(-242, 184) /w:[ -1 2 8 1 ]
  //: supply0 g19 (w36) @(-413,87) /sn:0 /w:[ 0 ]
  and g32 (.I0(w56), .I1(zero), .Z(w63));   //: @(-360,36) /sn:0 /w:[ 1 0 1 ]
  //: supply0 g38 (w9) @(-243,89) /sn:0 /w:[ 0 ]
  tran g6(.Z(w22), .I(IR[15:0]));   //: @(5,131) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g9(.Z(w37), .I(w22[15]));   //: @(92,272) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  //: supply1 g7 (w25) @(110,248) /sn:0 /w:[ 0 ]
  add g20 (.A(PC), .B(w49), .S(w46), .CI(w42), .CO(w48));   //: @(-208,358) /sn:0 /R:1 /w:[ 0 0 1 1 0 ]
  control g31 (.Op(Op), .Branch(w56), .RegWrite(WEN), .ALUSrc(w61), .ALUOp(w60), .MemWrite(w7), .MemToReg(w58), .MemRead(w57), .RegDest(w50));   //: @(-32, -94) /sz:(111, 110) /sn:0 /p:[ Bi0>1 Lo0<0 Ro0<0 Ro1<0 Ro2<0 Ro3<1 Ro4<0 Ro5<0 Ro6<0 ]
  //: supply1 g15 (w5) @(-147,54) /sn:0 /w:[ 0 ]
  //: joint g43 (reset) @(-51, 49) /w:[ 1 2 -1 8 ]
  //: joint g17 (PC) @(-242, 124) /w:[ 4 -1 6 3 ]
  //: dip g25 (w44) @(-333,414) /sn:0 /R:1 /w:[ 0 ] /st:2
  //: joint g29 (SB) @(92, 102) /w:[ 1 -1 2 4 ]
  //: joint g42 (clk) @(-46, 183) /w:[ 4 10 3 -1 ]
  //: joint g14 (Z) @(535, 161) /w:[ 2 4 -1 1 ]
  concat g5 (.I0(Inst), .I1(w13), .I2(w28), .I3(SB), .I4(SA), .I5(Op), .Z(IR));   //: @(42,107) /sn:0 /R:2 /w:[ 0 1 0 3 1 0 3 ] /dr:1
  //: supply0 g44 (w0) @(-194,190) /sn:0 /w:[ 0 ]
  //: joint g36 (clk) @(154, 183) /w:[ 6 -1 5 8 ]
  lshift g21 (.I(w24), .Z(w49), .S(w44));   //: @(-268,342) /sn:0 /R:1 /w:[ 5 1 1 ]
  //: supply0 g24 (w42) @(-194,328) /sn:0 /w:[ 0 ]
  //: supply0 g41 (w11) @(-26,101) /sn:0 /w:[ 1 ]
  mux g23 (.I0(w1), .I1(w46), .S(w63), .Z(nextPC));   //: @(-342,124) /sn:0 /R:1 /w:[ 1 0 0 0 ]
  //: joint g40 (reset) @(-281, -33) /w:[ 3 -1 4 6 ]
  clock g35 (.Z(clk));   //: @(-355,-1) /sn:0 /w:[ 0 ] /omega:800 /phi:0 /duty:50
  reg32 g0 (.WD(WD), .SA(SA), .SB(SB), .ENA(w4), .ENB(w4), .WA(WA), .WEN(WEN), .CLR(reset), .CLK(clk), .DA(A), .DB(w20));   //: @(185, 83) /sz:(99, 113) /sn:0 /p:[ Ti0>1 Li0>0 Li1>0 Li2>0 Li3>5 Li4>1 Li5>1 Li6>0 Li7>7 Bo0<0 Bo1<3 ]
  //: comment g26 /dolink:0 /link:"" @(-269,415) /sn:0 /R:1
  //: /line:"branch addr"
  //: /end
  //: joint g22 (w24) @(227, 269) /w:[ 2 -1 1 4 ]
  //: switch reset (reset) @(-356,-33) /sn:0 /w:[ 5 ] /st:0
  //: joint g12 (w20) @(255, 210) /w:[ 1 2 -1 4 ]
  //: dip g18 (w6) @(-507,82) /sn:0 /w:[ 0 ] /st:4
  ALU_control g30 (.ALUOp(w60), .Inst(Inst), .ALUop(ALUOp));   //: @(205, 327) /sz:(89, 65) /sn:0 /p:[ Ti0>1 Li0>1 Ro0<0 ]
  //: comment g33 /dolink:0 /link:"" @(-455,29) /sn:0
  //: /line:"alu zero"
  //: /end

endmodule

module reg32(CLR, DB, DA, CLK, WEN, WD, ENA, WA, ENB, SB, SA);
//: interface  /sz:(99, 111) /bd:[ Ti0>WD[31:0](47/99) Li0>SA[4:0](9/111) Li1>SB[4:0](19/111) Li2>ENA(37/111) Li3>ENB(47/111) Li4>WA[4:0](61/111) Li5>WEN(72/111) Li6>CLR(89/111) Li7>CLK(99/111) Bo0<DA[31:0](33/99) Bo1<DB[31:0](70/99) ]
input ENB;    //: /sn:0 {0}(56,99)(167,99)(167,106){1}
input [4:0] WA;    //: /sn:0 {0}(53,404)(65,404){1}
//: {2}(69,404)(82,404){3}
//: {4}(67,406)(67,436)(49,436)(49,451)(59,451){5}
input [31:0] WD;    //: /sn:0 {0}(518,185)(518,163)(294,163){1}
//: {2}(290,163)(140,163){3}
//: {4}(292,165)(292,184){5}
input [4:0] SB;    //: /sn:0 {0}(58,68)(83,68){1}
input CLR;    //: /sn:0 {0}(472,274)(451,274)(451,322)(235,322){1}
//: {2}(233,320)(233,273)(246,273){3}
//: {4}(231,322)(88,322){5}
input [4:0] SA;    //: /sn:0 {0}(74,-67)(102,-67){1}
input WEN;    //: /sn:0 {0}(69,485)(93,485){1}
output [31:0] DB;    //: /sn:0 /dp:1 {0}(550,298)(550,353){1}
//: {2}(552,355)(706,355){3}
//: {4}(548,355)(324,355)(324,297){5}
input CLK;    //: /sn:0 {0}(472,286)(461,286)(461,333)(241,333){1}
//: {2}(239,331)(239,285)(246,285){3}
//: {4}(237,333)(54,333){5}
output [31:0] DA;    //: /sn:0 /dp:1 {0}(280,297)(280,344)(504,344){1}
//: {2}(508,344)(705,344){3}
//: {4}(506,342)(506,298){5}
input ENA;    //: /sn:0 {0}(71,-42)(166,-42)(166,-33){1}
wire w6;    //: /sn:0 /dp:1 {0}(154,130)(137,130)(137,63)(89,63){1}
wire w7;    //: /sn:0 /dp:1 {0}(152,511)(120,511)(120,399)(88,399){1}
wire w4;    //: /sn:0 {0}(80,451)(86,451)(86,480)(93,480){1}
wire [3:0] w3;    //: /sn:0 {0}(246,194)(238,194)(238,-60){1}
//: {2}(240,-62)(467,-62)(467,195)(472,195){3}
//: {4}(236,-62)(108,-62){5}
wire w28;    //: /sn:0 {0}(181,521)(445,521)(445,260)(472,260){1}
wire w24;    //: /sn:0 {0}(183,140)(419,140)(419,233)(472,233){1}
wire w23;    //: /sn:0 {0}(183,120)(204,120)(204,232)(246,232){1}
wire w1;    //: /sn:0 /dp:1 {0}(153,-9)(144,-9)(144,-72)(108,-72){1}
wire w25;    //: /sn:0 {0}(114,483)(165,483)(165,487){1}
wire [3:0] w2;    //: /sn:0 {0}(89,73)(219,73){1}
//: {2}(223,73)(455,73)(455,207)(472,207){3}
//: {4}(221,75)(221,206)(246,206){5}
wire w12;    //: /sn:0 {0}(182,1)(431,1)(431,223)(472,223){1}
wire w27;    //: /sn:0 {0}(181,501)(227,501)(227,259)(246,259){1}
wire [3:0] w5;    //: /sn:0 {0}(88,409)(210,409){1}
//: {2}(214,409)(433,409)(433,250)(472,250){3}
//: {4}(212,407)(212,249)(246,249){5}
wire w9;    //: /sn:0 {0}(182,-19)(211,-19)(211,222)(246,222){1}
//: enddecls

  //: input g8 (CLR) @(86,322) /sn:0 /w:[ 5 ]
  //: joint g4 (DA) @(506, 344) /w:[ 2 4 1 -1 ]
  concat g13 (.I0(w3), .I1(w1), .Z(SA));   //: @(103,-67) /sn:0 /R:2 /w:[ 5 1 1 ] /dr:1
  //: output g3 (DB) @(703,355) /sn:0 /w:[ 3 ]
  //: output g2 (DA) @(702,344) /sn:0 /w:[ 3 ]
  reg16 g1 (.WD(WD), .SA(w3), .SB(w2), .ENA(w12), .ENB(w24), .WA(w5), .WEN(w28), .CLR(CLR), .CLK(CLK), .DA(DA), .DB(DB));   //: @(473, 186) /sz:(103, 111) /sn:0 /p:[ Ti0>0 Li0>3 Li1>3 Li2>1 Li3>1 Li4>3 Li5>1 Li6>0 Li7>0 Bo0<5 Bo1<0 ]
  demux g16 (.I(w1), .E(ENA), .Z0(w9), .Z1(w12));   //: @(166,-9) /sn:0 /R:1 /w:[ 0 1 0 0 ]
  //: joint g11 (CLK) @(239, 333) /w:[ 1 2 4 -1 ]
  and g28 (.I0(w4), .I1(WEN), .Z(w25));   //: @(104,483) /sn:0 /w:[ 1 1 0 ]
  //: input g10 (CLK) @(52,333) /sn:0 /w:[ 5 ]
  //: joint g32 (WA) @(67, 404) /w:[ 2 -1 1 4 ]
  //: input g27 (WEN) @(67,485) /sn:0 /w:[ 0 ]
  concat g19 (.I0(w2), .I1(w6), .Z(SB));   //: @(84,68) /sn:0 /R:2 /w:[ 0 1 1 ] /dr:1
  //: input g6 (WD) @(138,163) /sn:0 /w:[ 3 ]
  //: joint g9 (CLR) @(233, 322) /w:[ 1 2 4 -1 ]
  //: joint g7 (WD) @(292, 163) /w:[ 1 -1 2 4 ]
  or g31 (.I0(WA), .Z(w4));   //: @(70,451) /sn:0 /w:[ 5 0 ]
  //: input g15 (ENA) @(69,-42) /sn:0 /w:[ 0 ]
  //: joint g20 (w5) @(212, 409) /w:[ 2 4 1 -1 ]
  demux g29 (.I(w7), .E(w25), .Z0(w27), .Z1(w28));   //: @(165,511) /sn:0 /R:1 /w:[ 0 1 0 0 ]
  concat g25 (.I0(w5), .I1(w7), .Z(WA));   //: @(83,404) /sn:0 /R:2 /w:[ 0 1 3 ] /dr:1
  //: joint g17 (w2) @(221, 73) /w:[ 2 -1 1 4 ]
  //: joint g5 (DB) @(550, 355) /w:[ 2 1 4 -1 ]
  //: joint g14 (w3) @(238, -62) /w:[ 2 -1 4 1 ]
  //: input g24 (WA) @(51,404) /sn:0 /w:[ 0 ]
  demux g21 (.I(w6), .E(ENB), .Z0(w23), .Z1(w24));   //: @(167,130) /sn:0 /R:1 /w:[ 0 1 0 0 ]
  //: input g22 (ENB) @(54,99) /sn:0 /w:[ 0 ]
  reg16 g0 (.WD(WD), .SA(w3), .SB(w2), .ENA(w9), .ENB(w23), .WA(w5), .WEN(w27), .CLR(CLR), .CLK(CLK), .DA(DA), .DB(DB));   //: @(247, 185) /sz:(103, 111) /sn:0 /p:[ Ti0>5 Li0>0 Li1>5 Li2>1 Li3>1 Li4>5 Li5>1 Li6>3 Li7>3 Bo0<0 Bo1<5 ]
  //: input g18 (SB) @(56,68) /sn:0 /w:[ 0 ]
  //: input g12 (SA) @(72,-67) /sn:0 /w:[ 0 ]
  //: comment g33 /dolink:0 /link:"" @(5,524) /sn:0
  //: /line:"no writing to $0"
  //: /end

endmodule

module ALU_control(ALUop, Inst, ALUOp);
//: interface  /sz:(89, 65) /bd:[ Ti0>ALUOp[1:0](34/89) Li0>Inst[5:0](48/65) Ro0<ALUop[2:0](14/65) ]
output [2:0] ALUop;    //: /sn:0 /dp:1 {0}(419,208)(461,208){1}
input [5:0] Inst;    //: /sn:0 {0}(103,180)(122,180)(122,193){1}
//: {2}(122,194)(122,210){3}
//: {4}(122,211)(122,228){5}
//: {6}(122,229)(122,247){7}
//: {8}(122,248)(122,286){9}
input [1:0] ALUOp;    //: /sn:0 {0}(240,78)(258,78)(258,99){1}
//: {2}(258,100)(258,127){3}
//: {4}(258,128)(258,147){5}
wire w6;    //: /sn:0 {0}(400,169)(403,169)(403,198)(413,198){1}
wire w7;    //: /sn:0 {0}(126,248)(274,248){1}
wire w14;    //: /sn:0 {0}(353,244)(403,244)(403,218)(413,218){1}
wire w4;    //: /sn:0 {0}(262,100)(305,100)(305,166)(379,166){1}
wire w0;    //: /sn:0 {0}(332,241)(312,241)(312,212){1}
//: {2}(314,210)(338,210){3}
//: {4}(312,208)(312,174){5}
//: {6}(314,172)(337,172){7}
//: {8}(312,170)(312,128)(262,128){9}
wire w1;    //: /sn:0 {0}(126,194)(264,194)(264,243)(274,243){1}
wire w11;    //: /sn:0 {0}(295,246)(332,246){1}
wire w2;    //: /sn:0 /dp:1 {0}(337,177)(142,177)(142,211)(126,211){1}
wire w12;    //: /sn:0 {0}(359,208)(413,208){1}
wire w5;    //: /sn:0 {0}(338,205)(178,205)(178,229)(126,229){1}
wire w9;    //: /sn:0 {0}(358,175)(376,175)(376,171)(379,171){1}
//: enddecls

  or g4 (.I0(w1), .I1(w7), .Z(w11));   //: @(285,246) /sn:0 /w:[ 1 1 0 ]
  or g8 (.I0(!w5), .I1(!w0), .Z(w12));   //: @(349,208) /sn:0 /w:[ 0 3 0 ]
  //: output g3 (ALUop) @(458,208) /sn:0 /w:[ 1 ]
  or g13 (.I0(w4), .I1(w9), .Z(w6));   //: @(390,169) /sn:0 /w:[ 1 1 0 ]
  concat g2 (.I0(w14), .I1(w12), .I2(w6), .Z(ALUop));   //: @(418,208) /sn:0 /w:[ 1 1 1 0 ] /dr:0
  //: input g1 (Inst) @(101,180) /sn:0 /w:[ 0 ]
  tran g11(.Z(w4), .I(ALUOp[0]));   //: @(256,100) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: joint g10 (w0) @(312, 210) /w:[ 2 4 -1 1 ]
  tran g6(.Z(w5), .I(Inst[2]));   //: @(120,229) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  tran g9(.Z(w2), .I(Inst[1]));   //: @(120,211) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  and g7 (.I0(w0), .I1(w11), .Z(w14));   //: @(343,244) /sn:0 /w:[ 0 1 0 ]
  tran g15(.Z(w7), .I(Inst[3]));   //: @(120,248) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  and g17 (.I0(w0), .I1(w2), .Z(w9));   //: @(348,175) /sn:0 /w:[ 7 0 0 ]
  tran g5(.Z(w0), .I(ALUOp[1]));   //: @(256,128) /sn:0 /R:2 /w:[ 9 4 3 ] /ss:1
  tran g14(.Z(w1), .I(Inst[0]));   //: @(120,194) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: input g0 (ALUOp) @(238,78) /sn:0 /w:[ 0 ]
  //: comment g12 /dolink:0 /link:"" @(297,316) /sn:0
  //: /line:"1=!F2 or !Op1 or Op0"
  //: /end
  //: joint g18 (w0) @(312, 172) /w:[ 6 8 -1 5 ]

endmodule

module reg16(DA, ENA, SA, WD, DB, ENB, CLR, SB, WEN, CLK, WA);
//: interface  /sz:(103, 111) /bd:[ Ti0>WD[31:0](45/103) Li0>CLK(100/111) Li1>CLR(88/111) Li2>WEN(74/111) Li3>WA[3:0](64/111) Li4>ENB(47/111) Li5>ENA(37/111) Li6>SB[3:0](21/111) Li7>SA[3:0](9/111) Bo0<DB[31:0](77/103) Bo1<DA[31:0](33/103) ]
input ENB;    //: /sn:0 {0}(-22,52)(26,52)(26,56){1}
input [3:0] WA;    //: /sn:0 {0}(4,384)(37,384){1}
input [31:0] WD;    //: /sn:0 {0}(665,141)(665,124)(520,124){1}
//: {2}(516,124)(362,124){3}
//: {4}(358,124)(205,124){5}
//: {6}(201,124)(39,124){7}
//: {8}(203,126)(203,140){9}
//: {10}(360,126)(360,140){11}
//: {12}(518,126)(518,140){13}
input [3:0] SB;    //: /sn:0 {0}(-84,10)(-52,10){1}
input CLR;    //: /sn:0 {0}(615,233)(608,233)(608,291)(463,291){1}
//: {2}(461,289)(461,232)(468,232){3}
//: {4}(459,291)(305,291){5}
//: {6}(303,289)(303,232)(310,232){7}
//: {8}(301,291)(145,291){9}
//: {10}(143,289)(143,232)(153,232){11}
//: {12}(141,291)(41,291){13}
input [3:0] SA;    //: /sn:0 {0}(-57,-126)(-39,-126){1}
input WEN;    //: /sn:0 {0}(55,435)(87,435)(87,442){1}
output [31:0] DB;    //: /sn:0 /dp:1 {0}(232,251)(232,320)(387,320){1}
//: {2}(391,320)(545,320){3}
//: {4}(549,320)(692,320){5}
//: {6}(696,320)(768,320){7}
//: {8}(694,318)(694,252){9}
//: {10}(547,318)(547,251){11}
//: {12}(389,318)(389,251){13}
input CLK;    //: /sn:0 {0}(615,243)(612,243)(612,309)(467,309){1}
//: {2}(465,307)(465,242)(468,242){3}
//: {4}(463,309)(310,309){5}
//: {6}(308,307)(308,242)(310,242){7}
//: {8}(306,309)(151,309){9}
//: {10}(149,307)(149,242)(153,242){11}
//: {12}(147,309)(41,309){13}
output [31:0] DA;    //: /sn:0 /dp:1 {0}(184,251)(184,282)(339,282){1}
//: {2}(343,282)(497,282){3}
//: {4}(501,282)(644,282){5}
//: {6}(648,282)(767,282){7}
//: {8}(646,280)(646,252){9}
//: {10}(499,280)(499,251){11}
//: {12}(341,280)(341,251){13}
input ENA;    //: /sn:0 {0}(-45,-100)(24,-100)(24,-93){1}
wire w6;    //: /sn:0 {0}(42,62)(114,62)(114,187)(153,187){1}
wire w14;    //: /sn:0 {0}(42,74)(272,74)(272,187)(310,187){1}
wire w16;    //: /sn:0 {0}(103,460)(299,460)(299,213)(310,213){1}
wire w4;    //: /sn:0 {0}(103,448)(138,448)(138,213)(153,213){1}
wire [1:0] w31;    //: /sn:0 /dp:1 {0}(11,-69)(-1,-69)(-1,-131)(-33,-131){1}
wire w23;    //: /sn:0 {0}(42,86)(427,86)(427,187)(468,187){1}
wire [1:0] w1;    //: /sn:0 /dp:1 {0}(74,466)(67,466)(67,379)(43,379){1}
wire w25;    //: /sn:0 {0}(42,98)(580,98)(580,188)(615,188){1}
wire [1:0] w40;    //: /sn:0 /dp:1 {0}(13,80)(-2,80)(-2,5)(-46,5){1}
wire w8;    //: /sn:0 {0}(40,-87)(124,-87)(124,176)(153,176){1}
wire w22;    //: /sn:0 {0}(103,472)(457,472)(457,213)(468,213){1}
wire [1:0] w2;    //: /sn:0 {0}(-46,15)(133,15){1}
//: {2}(137,15)(290,15){3}
//: {4}(294,15)(444,15){5}
//: {6}(448,15)(606,15)(606,163)(615,163){7}
//: {8}(446,17)(446,162)(468,162){9}
//: {10}(292,17)(292,162)(310,162){11}
//: {12}(135,17)(135,162)(153,162){13}
wire w12;    //: /sn:0 {0}(40,-51)(588,-51)(588,177)(615,177){1}
wire [1:0] w11;    //: /sn:0 /dp:1 {0}(43,389)(118,389){1}
//: {2}(122,389)(284,389){3}
//: {4}(288,389)(442,389){5}
//: {6}(446,389)(593,389)(593,203)(615,203){7}
//: {8}(444,387)(444,202)(468,202){9}
//: {10}(286,387)(286,202)(310,202){11}
//: {12}(120,387)(120,202)(153,202){13}
wire w10;    //: /sn:0 {0}(40,-63)(437,-63)(437,176)(468,176){1}
wire w27;    //: /sn:0 {0}(103,484)(602,484)(602,214)(615,214){1}
wire [1:0] w13;    //: /sn:0 {0}(468,150)(459,150)(459,-119){1}
//: {2}(461,-121)(611,-121)(611,151)(615,151){3}
//: {4}(457,-121)(305,-121){5}
//: {6}(301,-121)(149,-121){7}
//: {8}(145,-121)(-33,-121){9}
//: {10}(147,-119)(147,150)(153,150){11}
//: {12}(303,-119)(303,150)(310,150){13}
wire w9;    //: /sn:0 {0}(40,-75)(283,-75)(283,176)(310,176){1}
//: enddecls

  //: output g8 (DA) @(764,282) /sn:0 /w:[ 7 ]
  reg4 g4 (.WD(WD), .SA(w13), .SB(w2), .ENA(w12), .ENB(w25), .WA(w11), .WEN(w27), .CLR(CLR), .CLK(CLK), .DA(DA), .DB(DB));   //: @(616, 142) /sz:(102, 109) /sn:0 /p:[ Ti0>0 Li0>3 Li1>7 Li2>1 Li3>1 Li4>7 Li5>1 Li6>0 Li7>0 Bo0<9 Bo1<9 ]
  //: input g13 (ENA) @(-47,-100) /sn:0 /w:[ 0 ]
  //: input g34 (SA) @(-59,-126) /sn:0 /w:[ 0 ]
  reg4 g3 (.WD(WD), .SA(w13), .SB(w2), .ENA(w10), .ENB(w23), .WA(w11), .WEN(w22), .CLR(CLR), .CLK(CLK), .DA(DA), .DB(DB));   //: @(469, 141) /sz:(102, 109) /sn:0 /p:[ Ti0>13 Li0>0 Li1>9 Li2>1 Li3>1 Li4>9 Li5>1 Li6>3 Li7>3 Bo0<11 Bo1<11 ]
  //: joint g37 (w13) @(147, -121) /w:[ 7 -1 8 10 ]
  reg4 g2 (.WD(WD), .SA(w13), .SB(w2), .ENA(w9), .ENB(w14), .WA(w11), .WEN(w16), .CLR(CLR), .CLK(CLK), .DA(DA), .DB(DB));   //: @(311, 141) /sz:(102, 109) /sn:0 /p:[ Ti0>11 Li0>13 Li1>11 Li2>1 Li3>1 Li4>11 Li5>1 Li6>7 Li7>7 Bo0<13 Bo1<13 ]
  //: input g1 (WD) @(37,124) /sn:0 /w:[ 7 ]
  //: output g16 (DB) @(765,320) /sn:0 /w:[ 7 ]
  //: joint g11 (DA) @(499, 282) /w:[ 4 10 3 -1 ]
  //: joint g10 (DB) @(694, 320) /w:[ 6 8 5 -1 ]
  concat g28 (.I0(w11), .I1(w1), .Z(WA));   //: @(38,384) /sn:0 /R:2 /w:[ 0 1 1 ] /dr:1
  demux g32 (.I(w1), .E(WEN), .Z0(w4), .Z1(w16), .Z2(w22), .Z3(w27));   //: @(87,466) /sn:0 /R:1 /w:[ 0 1 0 0 0 0 ]
  //: joint g27 (CLK) @(465, 309) /w:[ 1 2 4 -1 ]
  //: joint g19 (DB) @(389, 320) /w:[ 2 12 1 -1 ]
  //: input g38 (ENB) @(-24,52) /sn:0 /w:[ 0 ]
  //: joint g6 (WD) @(360, 124) /w:[ 3 -1 4 10 ]
  //: joint g9 (DA) @(646, 282) /w:[ 6 8 5 -1 ]
  //: joint g7 (WD) @(518, 124) /w:[ 1 -1 2 12 ]
  //: input g20 (CLR) @(39,291) /sn:0 /w:[ 13 ]
  //: joint g15 (w11) @(286, 389) /w:[ 4 10 3 -1 ]
  //: joint g31 (w11) @(120, 389) /w:[ 2 12 1 -1 ]
  //: input g39 (SB) @(-86,10) /sn:0 /w:[ 0 ]
  //: joint g43 (w2) @(446, 15) /w:[ 6 -1 5 8 ]
  //: input g29 (WEN) @(53,435) /sn:0 /w:[ 0 ]
  //: joint g25 (CLK) @(149, 309) /w:[ 9 10 12 -1 ]
  //: joint g17 (w13) @(459, -121) /w:[ 2 -1 4 1 ]
  //: joint g42 (w2) @(292, 15) /w:[ 4 -1 3 10 ]
  demux g14 (.I(w31), .E(ENA), .Z0(w8), .Z1(w9), .Z2(w10), .Z3(w12));   //: @(24,-69) /sn:0 /R:1 /w:[ 0 1 0 0 0 0 ]
  //: joint g5 (WD) @(203, 124) /w:[ 5 -1 6 8 ]
  //: joint g44 (w11) @(444, 389) /w:[ 6 8 5 -1 ]
  //: input g24 (CLK) @(39,309) /sn:0 /w:[ 13 ]
  //: joint g21 (CLR) @(143, 291) /w:[ 9 10 12 -1 ]
  //: joint g36 (w13) @(303, -121) /w:[ 5 -1 6 12 ]
  //: joint g23 (CLR) @(461, 291) /w:[ 1 2 4 -1 ]
  //: joint g41 (w2) @(135, 15) /w:[ 2 -1 1 12 ]
  concat g40 (.I0(w2), .I1(w40), .Z(SB));   //: @(-51,10) /sn:0 /R:2 /w:[ 0 1 1 ] /dr:1
  concat g35 (.I0(w13), .I1(w31), .Z(SA));   //: @(-38,-126) /sn:0 /R:2 /w:[ 9 1 1 ] /dr:1
  //: joint g26 (CLK) @(308, 309) /w:[ 5 6 8 -1 ]
  //: joint g22 (CLR) @(303, 291) /w:[ 5 6 8 -1 ]
  reg4 g0 (.WD(WD), .SA(w13), .SB(w2), .ENA(w8), .ENB(w6), .WA(w11), .WEN(w4), .CLR(CLR), .CLK(CLK), .DA(DA), .DB(DB));   //: @(154, 141) /sz:(102, 109) /sn:0 /p:[ Ti0>9 Li0>11 Li1>13 Li2>1 Li3>1 Li4>13 Li5>1 Li6>11 Li7>11 Bo0<0 Bo1<0 ]
  //: joint g18 (DB) @(547, 320) /w:[ 4 10 3 -1 ]
  //: joint g12 (DA) @(341, 282) /w:[ 2 12 1 -1 ]
  demux g33 (.I(w40), .E(ENB), .Z0(w6), .Z1(w14), .Z2(w23), .Z3(w25));   //: @(26,80) /sn:0 /R:1 /w:[ 0 1 0 0 0 0 ]
  //: input g30 (WA) @(2,384) /sn:0 /w:[ 0 ]

endmodule
